LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY clkdiv IS
PORT(CLK:IN STD_LOGIC;Q:OUT STD_LOGIC);
END clkdiv;
ARCHITECTURE BEHAV OF clkdiv IS
BEGIN 
PROCESS(CLK)
VARIABLE TIME:INTEGER RANGE 0 TO 50000000;
BEGIN
	IF RISING_EDGE(CLK) THEN
		TIME:=TIME+1;
		IF TIME=25000000 THEN
				Q<='1';
		ELSIF TIME=50000000 THEN
			Q<='0';
			TIME:=0;
		END IF;
	END IF;
END PROCESS;
END BEHAV;